module tpu_top#(
	parameter ARRAY_SIZE = 256,
	parameter SRAM_DATA_WIDTH = 32,
	parameter DATA_WIDTH = 8,
	parameter OUTPUT_DATA_WIDTH = 16
)
(
	input clk,
	input srstn,
	input tpu_start,

	//input data for (data, weight) from eight SRAM
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w0,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w1,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w2,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w3,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w4,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w5,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w6,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w7,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w8,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w9,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w10,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w11,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w12,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w13,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w14,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w15,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w16,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w17,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w18,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w19,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w20,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w21,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w22,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w23,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w24,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w25,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w26,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w27,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w28,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w29,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w30,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w31,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w32,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w33,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w34,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w35,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w36,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w37,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w38,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w39,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w40,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w41,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w42,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w43,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w44,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w45,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w46,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w47,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w48,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w49,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w50,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w51,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w52,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w53,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w54,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w55,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w56,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w57,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w58,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w59,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w60,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w61,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w62,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_w63,
	
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d0,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d1,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d2,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d3,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d4,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d5,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d6,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d7,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d8,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d9,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d10,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d11,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d12,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d13,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d14,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d15,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d16,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d17,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d18,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d19,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d20,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d21,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d22,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d23,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d24,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d25,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d26,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d27,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d28,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d29,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d30,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d31,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d32,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d33,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d34,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d35,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d36,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d37,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d38,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d39,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d40,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d41,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d42,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d43,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d44,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d45,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d46,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d47,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d48,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d49,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d50,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d51,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d52,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d53,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d54,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d55,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d56,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d57,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d58,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d59,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d60,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d61,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d62,
	input [SRAM_DATA_WIDTH-1:0] sram_rdata_d63,

	//output addr for (data, weight) from eight SRAM
	output [9:0] sram_raddr_w0,
	output [9:0] sram_raddr_w1,
	output [9:0] sram_raddr_w2,
	output [9:0] sram_raddr_w3,
	output [9:0] sram_raddr_w4,
	output [9:0] sram_raddr_w5,
	output [9:0] sram_raddr_w6,
	output [9:0] sram_raddr_w7,
	output [9:0] sram_raddr_w8,
	output [9:0] sram_raddr_w9,
	output [9:0] sram_raddr_w10,
	output [9:0] sram_raddr_w11,
	output [9:0] sram_raddr_w12,
	output [9:0] sram_raddr_w13,
	output [9:0] sram_raddr_w14,
	output [9:0] sram_raddr_w15,
	output [9:0] sram_raddr_w16,
	output [9:0] sram_raddr_w17,
	output [9:0] sram_raddr_w18,
	output [9:0] sram_raddr_w19,
	output [9:0] sram_raddr_w20,
	output [9:0] sram_raddr_w21,
	output [9:0] sram_raddr_w22,
	output [9:0] sram_raddr_w23,
	output [9:0] sram_raddr_w24,
	output [9:0] sram_raddr_w25,
	output [9:0] sram_raddr_w26,
	output [9:0] sram_raddr_w27,
	output [9:0] sram_raddr_w28,
	output [9:0] sram_raddr_w29,
	output [9:0] sram_raddr_w30,
	output [9:0] sram_raddr_w31,
	output [9:0] sram_raddr_w32,
	output [9:0] sram_raddr_w33,
	output [9:0] sram_raddr_w34,
	output [9:0] sram_raddr_w35,
	output [9:0] sram_raddr_w36,
	output [9:0] sram_raddr_w37,
	output [9:0] sram_raddr_w38,
	output [9:0] sram_raddr_w39,
	output [9:0] sram_raddr_w40,
	output [9:0] sram_raddr_w41,
	output [9:0] sram_raddr_w42,
	output [9:0] sram_raddr_w43,
	output [9:0] sram_raddr_w44,
	output [9:0] sram_raddr_w45,
	output [9:0] sram_raddr_w46,
	output [9:0] sram_raddr_w47,
	output [9:0] sram_raddr_w48,
	output [9:0] sram_raddr_w49,
	output [9:0] sram_raddr_w50,
	output [9:0] sram_raddr_w51,
	output [9:0] sram_raddr_w52,
	output [9:0] sram_raddr_w53,
	output [9:0] sram_raddr_w54,
	output [9:0] sram_raddr_w55,
	output [9:0] sram_raddr_w56,
	output [9:0] sram_raddr_w57,
	output [9:0] sram_raddr_w58,
	output [9:0] sram_raddr_w59,
	output [9:0] sram_raddr_w60,
	output [9:0] sram_raddr_w61,
	output [9:0] sram_raddr_w62,
	output [9:0] sram_raddr_w63,

	output [9:0] sram_raddr_d0,
	output [9:0] sram_raddr_d1,
	output [9:0] sram_raddr_d2,
	output [9:0] sram_raddr_d3,
	output [9:0] sram_raddr_d4,
	output [9:0] sram_raddr_d5,
	output [9:0] sram_raddr_d6,
	output [9:0] sram_raddr_d7,
	output [9:0] sram_raddr_d8,
	output [9:0] sram_raddr_d9,
	output [9:0] sram_raddr_d10,
	output [9:0] sram_raddr_d11,
	output [9:0] sram_raddr_d12,
	output [9:0] sram_raddr_d13,
	output [9:0] sram_raddr_d14,
	output [9:0] sram_raddr_d15,
	output [9:0] sram_raddr_d16,
	output [9:0] sram_raddr_d17,
	output [9:0] sram_raddr_d18,
	output [9:0] sram_raddr_d19,
	output [9:0] sram_raddr_d20,
	output [9:0] sram_raddr_d21,
	output [9:0] sram_raddr_d22,
	output [9:0] sram_raddr_d23,
	output [9:0] sram_raddr_d24,
	output [9:0] sram_raddr_d25,
	output [9:0] sram_raddr_d26,
	output [9:0] sram_raddr_d27,
	output [9:0] sram_raddr_d28,
	output [9:0] sram_raddr_d29,
	output [9:0] sram_raddr_d30,
	output [9:0] sram_raddr_d31,
	output [9:0] sram_raddr_d32,
	output [9:0] sram_raddr_d33,
	output [9:0] sram_raddr_d34,
	output [9:0] sram_raddr_d35,
	output [9:0] sram_raddr_d36,
	output [9:0] sram_raddr_d37,
	output [9:0] sram_raddr_d38,
	output [9:0] sram_raddr_d39,
	output [9:0] sram_raddr_d40,
	output [9:0] sram_raddr_d41,
	output [9:0] sram_raddr_d42,
	output [9:0] sram_raddr_d43,
	output [9:0] sram_raddr_d44,
	output [9:0] sram_raddr_d45,
	output [9:0] sram_raddr_d46,
	output [9:0] sram_raddr_d47,
	output [9:0] sram_raddr_d48,
	output [9:0] sram_raddr_d49,
	output [9:0] sram_raddr_d50,
	output [9:0] sram_raddr_d51,
	output [9:0] sram_raddr_d52,
	output [9:0] sram_raddr_d53,
	output [9:0] sram_raddr_d54,
	output [9:0] sram_raddr_d55,
	output [9:0] sram_raddr_d56,
	output [9:0] sram_raddr_d57,
	output [9:0] sram_raddr_d58,
	output [9:0] sram_raddr_d59,
	output [9:0] sram_raddr_d60,
	output [9:0] sram_raddr_d61,
	output [9:0] sram_raddr_d62,
	output [9:0] sram_raddr_d63,
	
	//write to three SRAN for comparison
	output sram_write_enable_a0,
	output [ARRAY_SIZE*OUTPUT_DATA_WIDTH-1:0] sram_wdata_a,
	output [5:0] sram_waddr_a,

	output sram_write_enable_b0,
	output [ARRAY_SIZE*OUTPUT_DATA_WIDTH-1:0] sram_wdata_b,
	output [5:0] sram_waddr_b,

	output sram_write_enable_c0,
	output [ARRAY_SIZE*OUTPUT_DATA_WIDTH-1:0] sram_wdata_c,
	output [5:0] sram_waddr_c,
	
	output tpu_done
);
localparam ORI_WIDTH = DATA_WIDTH+DATA_WIDTH+5;

//----addr_sel parameter----
wire [6:0] addr_serial_num;

//----quantized parameter----
wire signed [ARRAY_SIZE*ORI_WIDTH-1:0] ori_data;
wire signed [ARRAY_SIZE*OUTPUT_DATA_WIDTH-1:0] quantized_data;

//-----systolic parameter----
wire alu_start;
wire [8:0] cycle_num;
wire [5:0] matrix_index;

//----ststolic_controll parameter---
wire sram_write_enable;
wire [1:0] data_set;

//----write_out parameter----
// nothing XD



//----addr_sel module----
addr_sel addr_sel 
(
	//input
	.clk(clk),
	.addr_serial_num(addr_serial_num),	

	//output
	.sram_raddr_w0(sram_raddr_w0),
	.sram_raddr_w1(sram_raddr_w1),
	.sram_raddr_w2(sram_raddr_w2),
	.sram_raddr_w3(sram_raddr_w3),
	.sram_raddr_w4(sram_raddr_w4),
	.sram_raddr_w5(sram_raddr_w5),
	.sram_raddr_w6(sram_raddr_w6),
	.sram_raddr_w7(sram_raddr_w7),
	.sram_raddr_w8(sram_raddr_w8),
	.sram_raddr_w9(sram_raddr_w9),
	.sram_raddr_w10(sram_raddr_w10),
	.sram_raddr_w11(sram_raddr_w11),
	.sram_raddr_w12(sram_raddr_w12),
	.sram_raddr_w13(sram_raddr_w13),
	.sram_raddr_w14(sram_raddr_w14),
	.sram_raddr_w15(sram_raddr_w15),
	.sram_raddr_w16(sram_raddr_w16),
	.sram_raddr_w17(sram_raddr_w17),
	.sram_raddr_w18(sram_raddr_w18),
	.sram_raddr_w19(sram_raddr_w19),
	.sram_raddr_w20(sram_raddr_w20),
	.sram_raddr_w21(sram_raddr_w21),
	.sram_raddr_w22(sram_raddr_w22),
	.sram_raddr_w23(sram_raddr_w23),
	.sram_raddr_w24(sram_raddr_w24),
	.sram_raddr_w25(sram_raddr_w25),
	.sram_raddr_w26(sram_raddr_w26),
	.sram_raddr_w27(sram_raddr_w27),
	.sram_raddr_w28(sram_raddr_w28),
	.sram_raddr_w29(sram_raddr_w29),
	.sram_raddr_w30(sram_raddr_w30),
	.sram_raddr_w31(sram_raddr_w31),
	.sram_raddr_w32(sram_raddr_w32),
	.sram_raddr_w33(sram_raddr_w33),
	.sram_raddr_w34(sram_raddr_w34),
	.sram_raddr_w35(sram_raddr_w35),
	.sram_raddr_w36(sram_raddr_w36),
	.sram_raddr_w37(sram_raddr_w37),
	.sram_raddr_w38(sram_raddr_w38),
	.sram_raddr_w39(sram_raddr_w39),
	.sram_raddr_w40(sram_raddr_w40),
	.sram_raddr_w41(sram_raddr_w41),
	.sram_raddr_w42(sram_raddr_w42),
	.sram_raddr_w43(sram_raddr_w43),
	.sram_raddr_w44(sram_raddr_w44),
	.sram_raddr_w45(sram_raddr_w45),
	.sram_raddr_w46(sram_raddr_w46),
	.sram_raddr_w47(sram_raddr_w47),
	.sram_raddr_w48(sram_raddr_w48),
	.sram_raddr_w49(sram_raddr_w49),
	.sram_raddr_w50(sram_raddr_w50),
	.sram_raddr_w51(sram_raddr_w51),
	.sram_raddr_w52(sram_raddr_w52),
	.sram_raddr_w53(sram_raddr_w53),
	.sram_raddr_w54(sram_raddr_w54),
	.sram_raddr_w55(sram_raddr_w55),
	.sram_raddr_w56(sram_raddr_w56),
	.sram_raddr_w57(sram_raddr_w57),
	.sram_raddr_w58(sram_raddr_w58),
	.sram_raddr_w59(sram_raddr_w59),
	.sram_raddr_w60(sram_raddr_w60),
	.sram_raddr_w61(sram_raddr_w61),
	.sram_raddr_w62(sram_raddr_w62),
	.sram_raddr_w63(sram_raddr_w63),

	.sram_raddr_d0(sram_raddr_d0),
	.sram_raddr_d1(sram_raddr_d1),
	.sram_raddr_d2(sram_raddr_d2),
	.sram_raddr_d3(sram_raddr_d3),
	.sram_raddr_d4(sram_raddr_d4),
	.sram_raddr_d5(sram_raddr_d5),
	.sram_raddr_d6(sram_raddr_d6),
	.sram_raddr_d7(sram_raddr_d7),
	.sram_raddr_d8(sram_raddr_d8),
	.sram_raddr_d9(sram_raddr_d9),
	.sram_raddr_d10(sram_raddr_d10),
	.sram_raddr_d11(sram_raddr_d11),
	.sram_raddr_d12(sram_raddr_d12),
	.sram_raddr_d13(sram_raddr_d13),
	.sram_raddr_d14(sram_raddr_d14),
	.sram_raddr_d15(sram_raddr_d15),
	.sram_raddr_d16(sram_raddr_d16),
	.sram_raddr_d17(sram_raddr_d17),
	.sram_raddr_d18(sram_raddr_d18),
	.sram_raddr_d19(sram_raddr_d19),
	.sram_raddr_d20(sram_raddr_d20),
	.sram_raddr_d21(sram_raddr_d21),
	.sram_raddr_d22(sram_raddr_d22),
	.sram_raddr_d23(sram_raddr_d23),
	.sram_raddr_d24(sram_raddr_d24),
	.sram_raddr_d25(sram_raddr_d25),
	.sram_raddr_d26(sram_raddr_d26),
	.sram_raddr_d27(sram_raddr_d27),
	.sram_raddr_d28(sram_raddr_d28),
	.sram_raddr_d29(sram_raddr_d29),
	.sram_raddr_d30(sram_raddr_d30),
	.sram_raddr_d31(sram_raddr_d31),
	.sram_raddr_d32(sram_raddr_d32),
	.sram_raddr_d33(sram_raddr_d33),
	.sram_raddr_d34(sram_raddr_d34),
	.sram_raddr_d35(sram_raddr_d35),
	.sram_raddr_d36(sram_raddr_d36),
	.sram_raddr_d37(sram_raddr_d37),
	.sram_raddr_d38(sram_raddr_d38),
	.sram_raddr_d39(sram_raddr_d39),
	.sram_raddr_d40(sram_raddr_d40),
	.sram_raddr_d41(sram_raddr_d41),
	.sram_raddr_d42(sram_raddr_d42),
	.sram_raddr_d43(sram_raddr_d43),
	.sram_raddr_d44(sram_raddr_d44),
	.sram_raddr_d45(sram_raddr_d45),
	.sram_raddr_d46(sram_raddr_d46),
	.sram_raddr_d47(sram_raddr_d47),
	.sram_raddr_d48(sram_raddr_d48),
	.sram_raddr_d49(sram_raddr_d49),
	.sram_raddr_d50(sram_raddr_d50),
	.sram_raddr_d51(sram_raddr_d51),
	.sram_raddr_d52(sram_raddr_d52),
	.sram_raddr_d53(sram_raddr_d53),
	.sram_raddr_d54(sram_raddr_d54),
	.sram_raddr_d55(sram_raddr_d55),
	.sram_raddr_d56(sram_raddr_d56),
	.sram_raddr_d57(sram_raddr_d57),
	.sram_raddr_d58(sram_raddr_d58),
	.sram_raddr_d59(sram_raddr_d59),
	.sram_raddr_d60(sram_raddr_d60),
	.sram_raddr_d61(sram_raddr_d61),
	.sram_raddr_d62(sram_raddr_d62),
	.sram_raddr_d63(sram_raddr_d63)
);

//----quantize module----
quantize #(
	.ARRAY_SIZE(ARRAY_SIZE),
	.SRAM_DATA_WIDTH(SRAM_DATA_WIDTH),
	.DATA_WIDTH(DATA_WIDTH),
	.OUTPUT_DATA_WIDTH(OUTPUT_DATA_WIDTH)
) quantize
(
	//input
	.ori_data(ori_data),

	//output
	.quantized_data(quantized_data)	
);

//----systolic module----
systolic #(
	.ARRAY_SIZE(ARRAY_SIZE),
	.SRAM_DATA_WIDTH(SRAM_DATA_WIDTH),
	.DATA_WIDTH(DATA_WIDTH)
) systolic
(
	//input
	.clk(clk),
	.srstn(srstn),
	.alu_start(alu_start),
	.cycle_num(cycle_num),

	.sram_rdata_w0(sram_rdata_w0),
	.sram_rdata_w1(sram_rdata_w1),
	.sram_rdata_w2(sram_rdata_w2),
	.sram_rdata_w3(sram_rdata_w3),
	.sram_rdata_w4(sram_rdata_w4),
	.sram_rdata_w5(sram_rdata_w5),
	.sram_rdata_w6(sram_rdata_w6),
	.sram_rdata_w7(sram_rdata_w7),
	.sram_rdata_w8(sram_rdata_w8),
	.sram_rdata_w9(sram_rdata_w9),
	.sram_rdata_w10(sram_rdata_w10),
	.sram_rdata_w11(sram_rdata_w11),
	.sram_rdata_w12(sram_rdata_w12),
	.sram_rdata_w13(sram_rdata_w13),
	.sram_rdata_w14(sram_rdata_w14),
	.sram_rdata_w15(sram_rdata_w15),
	.sram_rdata_w16(sram_rdata_w16),
	.sram_rdata_w17(sram_rdata_w17),
	.sram_rdata_w18(sram_rdata_w18),
	.sram_rdata_w19(sram_rdata_w19),
	.sram_rdata_w20(sram_rdata_w20),
	.sram_rdata_w21(sram_rdata_w21),
	.sram_rdata_w22(sram_rdata_w22),
	.sram_rdata_w23(sram_rdata_w23),
	.sram_rdata_w24(sram_rdata_w24),
	.sram_rdata_w25(sram_rdata_w25),
	.sram_rdata_w26(sram_rdata_w26),
	.sram_rdata_w27(sram_rdata_w27),
	.sram_rdata_w28(sram_rdata_w28),
	.sram_rdata_w29(sram_rdata_w29),
	.sram_rdata_w30(sram_rdata_w30),
	.sram_rdata_w31(sram_rdata_w31),
	.sram_rdata_w32(sram_rdata_w32),
	.sram_rdata_w33(sram_rdata_w33),
	.sram_rdata_w34(sram_rdata_w34),
	.sram_rdata_w35(sram_rdata_w35),
	.sram_rdata_w36(sram_rdata_w36),
	.sram_rdata_w37(sram_rdata_w37),
	.sram_rdata_w38(sram_rdata_w38),
	.sram_rdata_w39(sram_rdata_w39),
	.sram_rdata_w40(sram_rdata_w40),
	.sram_rdata_w41(sram_rdata_w41),
	.sram_rdata_w42(sram_rdata_w42),
	.sram_rdata_w43(sram_rdata_w43),
	.sram_rdata_w44(sram_rdata_w44),
	.sram_rdata_w45(sram_rdata_w45),
	.sram_rdata_w46(sram_rdata_w46),
	.sram_rdata_w47(sram_rdata_w47),
	.sram_rdata_w48(sram_rdata_w48),
	.sram_rdata_w49(sram_rdata_w49),
	.sram_rdata_w50(sram_rdata_w50),
	.sram_rdata_w51(sram_rdata_w51),
	.sram_rdata_w52(sram_rdata_w52),
	.sram_rdata_w53(sram_rdata_w53),
	.sram_rdata_w54(sram_rdata_w54),
	.sram_rdata_w55(sram_rdata_w55),
	.sram_rdata_w56(sram_rdata_w56),
	.sram_rdata_w57(sram_rdata_w57),
	.sram_rdata_w58(sram_rdata_w58),
	.sram_rdata_w59(sram_rdata_w59),
	.sram_rdata_w60(sram_rdata_w60),
	.sram_rdata_w61(sram_rdata_w61),
	.sram_rdata_w62(sram_rdata_w62),
	.sram_rdata_w63(sram_rdata_w63),
		
	.sram_rdata_d0(sram_rdata_d0),
	.sram_rdata_d1(sram_rdata_d1),
	.sram_rdata_d2(sram_rdata_d2),
	.sram_rdata_d3(sram_rdata_d3),
	.sram_rdata_d4(sram_rdata_d4),
	.sram_rdata_d5(sram_rdata_d5),
	.sram_rdata_d6(sram_rdata_d6),
	.sram_rdata_d7(sram_rdata_d7),
	.sram_rdata_d8(sram_rdata_d8),
	.sram_rdata_d9(sram_rdata_d9),
	.sram_rdata_d10(sram_rdata_d10),
	.sram_rdata_d11(sram_rdata_d11),
	.sram_rdata_d12(sram_rdata_d12),
	.sram_rdata_d13(sram_rdata_d13),
	.sram_rdata_d14(sram_rdata_d14),
	.sram_rdata_d15(sram_rdata_d15),
	.sram_rdata_d16(sram_rdata_d16),
	.sram_rdata_d17(sram_rdata_d17),
	.sram_rdata_d18(sram_rdata_d18),
	.sram_rdata_d19(sram_rdata_d19),
	.sram_rdata_d20(sram_rdata_d20),
	.sram_rdata_d21(sram_rdata_d21),
	.sram_rdata_d22(sram_rdata_d22),
	.sram_rdata_d23(sram_rdata_d23),
	.sram_rdata_d24(sram_rdata_d24),
	.sram_rdata_d25(sram_rdata_d25),
	.sram_rdata_d26(sram_rdata_d26),
	.sram_rdata_d27(sram_rdata_d27),
	.sram_rdata_d28(sram_rdata_d28),
	.sram_rdata_d29(sram_rdata_d29),
	.sram_rdata_d30(sram_rdata_d30),
	.sram_rdata_d31(sram_rdata_d31),
	.sram_rdata_d32(sram_rdata_d32),
	.sram_rdata_d33(sram_rdata_d33),
	.sram_rdata_d34(sram_rdata_d34),
	.sram_rdata_d35(sram_rdata_d35),
	.sram_rdata_d36(sram_rdata_d36),
	.sram_rdata_d37(sram_rdata_d37),
	.sram_rdata_d38(sram_rdata_d38),
	.sram_rdata_d39(sram_rdata_d39),
	.sram_rdata_d40(sram_rdata_d40),
	.sram_rdata_d41(sram_rdata_d41),
	.sram_rdata_d42(sram_rdata_d42),
	.sram_rdata_d43(sram_rdata_d43),
	.sram_rdata_d44(sram_rdata_d44),
	.sram_rdata_d45(sram_rdata_d45),
	.sram_rdata_d46(sram_rdata_d46),
	.sram_rdata_d47(sram_rdata_d47),
	.sram_rdata_d48(sram_rdata_d48),
	.sram_rdata_d49(sram_rdata_d49),
	.sram_rdata_d50(sram_rdata_d50),
	.sram_rdata_d51(sram_rdata_d51),
	.sram_rdata_d52(sram_rdata_d52),
	.sram_rdata_d53(sram_rdata_d53),
	.sram_rdata_d54(sram_rdata_d54),
	.sram_rdata_d55(sram_rdata_d55),
	.sram_rdata_d56(sram_rdata_d56),
	.sram_rdata_d57(sram_rdata_d57),
	.sram_rdata_d58(sram_rdata_d58),
	.sram_rdata_d59(sram_rdata_d59),
	.sram_rdata_d60(sram_rdata_d60),
	.sram_rdata_d61(sram_rdata_d61),
	.sram_rdata_d62(sram_rdata_d62),
	.sram_rdata_d63(sram_rdata_d63),

	.matrix_index(matrix_index),
	
	//output
	.mul_outcome(ori_data)
);

//----systolic_controller module----
systolic_controll  #(
	.ARRAY_SIZE(ARRAY_SIZE)
) systolic_controll
(
	//input
	.clk(clk),
	.srstn(srstn),
	.tpu_start(tpu_start),

	//output
	.sram_write_enable(sram_write_enable),
	.addr_serial_num(addr_serial_num),
	.alu_start(alu_start),
	.cycle_num(cycle_num),
	.matrix_index(matrix_index),
	.data_set(data_set),
	.tpu_done(tpu_done)
);

//----write_out module----
write_out #(
	.ARRAY_SIZE(ARRAY_SIZE),
	.OUTPUT_DATA_WIDTH(OUTPUT_DATA_WIDTH)
) write_out
(
	//input
	.clk(clk), 
	.srstn(srstn),
	.sram_write_enable(sram_write_enable),
	.data_set(data_set),
	.matrix_index(matrix_index),
	.quantized_data(quantized_data),

	//output
	.sram_write_enable_a0(sram_write_enable_a0),
	.sram_wdata_a(sram_wdata_a),
	.sram_waddr_a(sram_waddr_a),

	.sram_write_enable_b0(sram_write_enable_b0),
	.sram_wdata_b(sram_wdata_b),
	.sram_waddr_b(sram_waddr_b),

	.sram_write_enable_c0(sram_write_enable_c0),
	.sram_wdata_c(sram_wdata_c),
	.sram_waddr_c(sram_waddr_c)
);

endmodule

